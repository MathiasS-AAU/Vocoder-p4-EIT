----------------------------------------------------------------------------------
-- Company:				AAU
-- Engineer: 			EIT4-415
-- Create Date:    	15/04/2020 
-- Design Name: 	 	Control Unit
-- Module Name:    	CU - control_unit - Behavioral 
-- Description:		The Finite State Machine controlling the data path and
--							memory, based on hardcoded instructions
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity control_unit is
end control_unit;

architecture Behavioral of control_unit is

begin


end Behavioral;

