----------------------------------------------------------------------------------
-- Company:				AAU
-- Engineer: 			EIT4-415
-- Create Date:    	15/04/2020 
-- Design Name: 	 	Arithmetic Logic Unit
-- Module Name:    	ALU - ALU - Behavioral
-- Description:		A signal from control unit will determine which operation
--							to execute
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ALU is
end ALU;

architecture Behavioral of ALU is

begin


end Behavioral;

