----------------------------------------------------------------------------------
-- Company:				AAU
-- Engineer: 			EIT4-415
-- Create Date:    	15/04/2020 
-- Design Name: 	 	Program Memory
-- Module Name:    	ROM - rom_32733x16_sync - Behavioral 
-- Description:		Read Only Memory (Don't overwrite the program!)
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity rom_32733x16_sync is
end rom_32733x16_sync;

architecture Behavioral of rom_32733x16_sync is

begin


end Behavioral;

